magic
tech sky130A
timestamp 1612933953
<< nwell >>
rect -120 195 150 335
<< nmos >>
rect 0 0 15 100
rect 40 0 55 100
<< pmos >>
rect 0 215 15 315
rect 65 215 80 315
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 100
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
<< pdiff >>
rect -50 300 0 315
rect -50 230 -35 300
rect -15 230 0 300
rect -50 215 0 230
rect 15 300 65 315
rect 15 230 30 300
rect 50 230 65 300
rect 15 215 65 230
rect 80 300 130 315
rect 80 230 95 300
rect 115 230 130 300
rect 80 215 130 230
<< ndiffc >>
rect -35 15 -15 85
rect 70 15 90 85
<< pdiffc >>
rect -35 230 -15 300
rect 30 230 50 300
rect 95 230 115 300
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 300 -50 315
rect -100 230 -85 300
rect -65 230 -50 300
rect -100 215 -50 230
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 230 -65 300
<< poly >>
rect 0 315 15 330
rect 65 315 80 330
rect 0 100 15 215
rect 65 130 80 215
rect 40 115 80 130
rect 40 100 55 115
rect 0 -15 15 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
rect 40 -80 55 0
rect 15 -90 55 -80
rect 15 -110 25 -90
rect 45 -110 55 -90
rect 15 -120 55 -110
<< polycont >>
rect -15 -45 5 -25
rect 25 -110 45 -90
<< locali >>
rect -95 300 -5 310
rect -95 230 -85 300
rect -65 230 -35 300
rect -15 230 -5 300
rect -95 220 -5 230
rect 20 300 60 310
rect 20 230 30 300
rect 50 230 60 300
rect 20 220 60 230
rect 85 300 125 310
rect 85 230 95 300
rect 115 230 125 300
rect 85 220 125 230
rect 40 95 60 220
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect 40 85 100 95
rect 40 75 70 85
rect -95 5 -5 15
rect 60 15 70 75
rect 90 15 100 85
rect 60 5 100 15
rect 80 -15 100 5
rect -120 -25 15 -15
rect -120 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 80 -35 150 -15
rect -25 -55 15 -45
rect -120 -90 55 -80
rect -120 -100 25 -90
rect 15 -110 25 -100
rect 45 -110 55 -90
rect 15 -120 55 -110
<< viali >>
rect -85 230 -65 300
rect -35 230 -15 300
rect 95 230 115 300
rect -85 15 -65 85
rect -35 15 -15 85
<< metal1 >>
rect -120 300 150 310
rect -120 230 -85 300
rect -65 230 -35 300
rect -15 230 95 300
rect 115 230 150 300
rect -120 220 150 230
rect -120 85 150 95
rect -120 15 -85 85
rect -65 15 -35 85
rect -15 15 150 85
rect -120 5 150 15
<< end >>
