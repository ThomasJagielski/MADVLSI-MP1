magic
tech sky130A
timestamp 1613052865
<< nwell >>
rect -120 235 85 475
<< nmos >>
rect 0 100 15 200
<< pmos >>
rect 0 255 15 455
<< ndiff >>
rect -50 185 0 200
rect -50 115 -35 185
rect -15 115 0 185
rect -50 100 0 115
rect 15 185 65 200
rect 15 115 30 185
rect 50 115 65 185
rect 15 100 65 115
<< pdiff >>
rect -50 440 0 455
rect -50 370 -35 440
rect -15 370 0 440
rect -50 340 0 370
rect -50 270 -35 340
rect -15 270 0 340
rect -50 255 0 270
rect 15 440 65 455
rect 15 370 30 440
rect 50 370 65 440
rect 15 340 65 370
rect 15 270 30 340
rect 50 270 65 340
rect 15 255 65 270
<< ndiffc >>
rect -35 115 -15 185
rect 30 115 50 185
<< pdiffc >>
rect -35 370 -15 440
rect -35 270 -15 340
rect 30 370 50 440
rect 30 270 50 340
<< psubdiff >>
rect -100 185 -50 200
rect -100 115 -85 185
rect -65 115 -50 185
rect -100 100 -50 115
<< nsubdiff >>
rect -100 440 -50 455
rect -100 370 -85 440
rect -65 370 -50 440
rect -100 340 -50 370
rect -100 270 -85 340
rect -65 270 -50 340
rect -100 255 -50 270
<< psubdiffcont >>
rect -85 115 -65 185
<< nsubdiffcont >>
rect -85 370 -65 440
rect -85 270 -65 340
<< poly >>
rect 0 455 15 470
rect 0 200 15 255
rect 0 -15 15 100
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
<< polycont >>
rect -15 -45 5 -25
<< locali >>
rect -95 440 -5 450
rect -95 370 -85 440
rect -65 370 -35 440
rect -15 370 -5 440
rect -95 340 -5 370
rect -95 270 -85 340
rect -65 270 -35 340
rect -15 270 -5 340
rect -95 260 -5 270
rect 20 440 60 450
rect 20 370 30 440
rect 50 370 60 440
rect 20 340 60 370
rect 20 270 30 340
rect 50 270 60 340
rect 20 260 60 270
rect 40 195 60 260
rect -95 185 -5 195
rect -95 115 -85 185
rect -65 115 -35 185
rect -15 115 -5 185
rect -95 105 -5 115
rect 20 185 60 195
rect 20 115 30 185
rect 50 115 60 185
rect 20 105 60 115
rect 40 -15 60 105
rect -120 -25 15 -15
rect -120 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 40 -35 85 -15
rect -25 -55 15 -45
<< viali >>
rect -85 370 -65 440
rect -35 370 -15 440
rect -85 270 -65 340
rect -35 270 -15 340
rect -85 115 -65 185
rect -35 115 -15 185
<< metal1 >>
rect -120 440 85 450
rect -120 370 -85 440
rect -65 370 -35 440
rect -15 370 85 440
rect -120 340 85 370
rect -120 270 -85 340
rect -65 270 -35 340
rect -15 270 85 340
rect -120 260 85 270
rect -120 185 85 195
rect -120 115 -85 185
rect -65 115 -35 185
rect -15 115 85 185
rect -120 5 85 115
<< labels >>
rlabel metal1 -120 100 -120 100 7 VN
port 4 w
rlabel locali 85 -25 85 -25 3 Y
port 2 e
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel metal1 -120 355 -120 355 7 VP
port 3 w
<< end >>
