magic
tech sky130A
timestamp 1612972315
<< nwell >>
rect -120 410 150 650
<< nmos >>
rect 25 60 40 260
rect 65 60 80 260
<< pmos >>
rect 0 430 15 630
rect 65 430 80 630
<< ndiff >>
rect -25 245 25 260
rect -25 175 -10 245
rect 10 175 25 245
rect -25 145 25 175
rect -25 75 -10 145
rect 10 75 25 145
rect -25 60 25 75
rect 40 60 65 260
rect 80 245 130 260
rect 80 175 95 245
rect 115 175 130 245
rect 80 145 130 175
rect 80 75 95 145
rect 115 75 130 145
rect 80 60 130 75
<< pdiff >>
rect -50 615 0 630
rect -50 545 -35 615
rect -15 545 0 615
rect -50 515 0 545
rect -50 445 -35 515
rect -15 445 0 515
rect -50 430 0 445
rect 15 615 65 630
rect 15 545 30 615
rect 50 545 65 615
rect 15 515 65 545
rect 15 445 30 515
rect 50 445 65 515
rect 15 430 65 445
rect 80 615 130 630
rect 80 545 95 615
rect 115 545 130 615
rect 80 515 130 545
rect 80 445 95 515
rect 115 445 130 515
rect 80 430 130 445
<< ndiffc >>
rect -10 175 10 245
rect -10 75 10 145
rect 95 175 115 245
rect 95 75 115 145
<< pdiffc >>
rect -35 545 -15 615
rect -35 445 -15 515
rect 30 545 50 615
rect 30 445 50 515
rect 95 545 115 615
rect 95 445 115 515
<< psubdiff >>
rect -75 245 -25 260
rect -75 175 -60 245
rect -40 175 -25 245
rect -75 145 -25 175
rect -75 75 -60 145
rect -40 75 -25 145
rect -75 60 -25 75
<< nsubdiff >>
rect -100 615 -50 630
rect -100 545 -85 615
rect -65 545 -50 615
rect -100 515 -50 545
rect -100 445 -85 515
rect -65 445 -50 515
rect -100 430 -50 445
<< psubdiffcont >>
rect -60 175 -40 245
rect -60 75 -40 145
<< nsubdiffcont >>
rect -85 545 -65 615
rect -85 445 -65 515
<< poly >>
rect 0 630 15 645
rect 65 630 80 645
rect 0 410 15 430
rect -25 400 15 410
rect -25 380 -15 400
rect 5 380 15 400
rect -25 370 15 380
rect 0 285 15 370
rect 65 350 80 430
rect 40 340 80 350
rect 40 320 50 340
rect 70 320 80 340
rect 40 310 80 320
rect 0 270 40 285
rect 25 260 40 270
rect 65 260 80 310
rect 25 45 40 60
rect 65 45 80 60
<< polycont >>
rect -15 380 5 400
rect 50 320 70 340
<< locali >>
rect -95 615 -5 625
rect -95 545 -85 615
rect -65 545 -35 615
rect -15 545 -5 615
rect -95 515 -5 545
rect -95 445 -85 515
rect -65 445 -35 515
rect -15 445 -5 515
rect -95 435 -5 445
rect 20 615 60 625
rect 20 545 30 615
rect 50 545 60 615
rect 20 515 60 545
rect 20 445 30 515
rect 50 445 60 515
rect 20 435 60 445
rect 85 615 125 625
rect 85 545 95 615
rect 115 545 125 615
rect 85 515 125 545
rect 85 445 95 515
rect 115 445 125 515
rect 85 435 125 445
rect 40 410 60 435
rect -120 400 15 410
rect -120 390 -15 400
rect -25 380 -15 390
rect 5 380 15 400
rect 40 390 150 410
rect -25 370 15 380
rect 40 340 80 350
rect 40 330 50 340
rect -120 320 50 330
rect 70 320 80 340
rect -120 310 80 320
rect 105 255 125 390
rect -70 245 20 255
rect -70 175 -60 245
rect -40 175 -10 245
rect 10 175 20 245
rect -70 145 20 175
rect -70 75 -60 145
rect -40 75 -10 145
rect 10 75 20 145
rect -70 65 20 75
rect 85 245 125 255
rect 85 175 95 245
rect 115 175 125 245
rect 85 145 125 175
rect 85 75 95 145
rect 115 75 125 145
rect 85 65 125 75
<< viali >>
rect -85 545 -65 615
rect -35 545 -15 615
rect -85 445 -65 515
rect -35 445 -15 515
rect 95 545 115 615
rect 95 445 115 515
rect -60 175 -40 245
rect -10 175 10 245
rect -60 75 -40 145
rect -10 75 10 145
<< metal1 >>
rect -120 615 150 625
rect -120 545 -85 615
rect -65 545 -35 615
rect -15 545 95 615
rect 115 545 150 615
rect -120 515 150 545
rect -120 445 -85 515
rect -65 445 -35 515
rect -15 445 95 515
rect 115 445 150 515
rect -120 435 150 445
rect -120 245 150 255
rect -120 175 -60 245
rect -40 175 -10 245
rect 10 175 150 245
rect -120 145 150 175
rect -120 75 -60 145
rect -40 75 -10 145
rect 10 75 150 145
rect -120 65 150 75
<< labels >>
rlabel locali -120 400 -120 400 7 A
port 1 w
rlabel locali -120 320 -120 320 7 B
port 2 w
rlabel locali 150 400 150 400 3 Y
port 3 e
rlabel metal1 -120 530 -120 530 7 VP
port 4 w
rlabel metal1 -120 160 -120 160 7 VN
port 5 w
<< end >>
